library verilog;
use verilog.vl_types.all;
entity qq_v is
end qq_v;
