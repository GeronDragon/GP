library verilog;
use verilog.vl_types.all;
entity test_v is
end test_v;
