library verilog;
use verilog.vl_types.all;
entity tt_v is
end tt_v;
